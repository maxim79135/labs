schp_inst : schp PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		enable	 => enable_sig,
		sclr	 => sclr_sig,
		q	 => q_sig
	);
