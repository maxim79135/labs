or5har_inst : or5har PORT MAP (
		data	 => data_sig,
		result	 => result_sig
	);
