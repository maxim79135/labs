sm2_inst : sm2 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		cout	 => cout_sig,
		result	 => result_sig
	);
