inector11_inst : inector11 PORT MAP (
		data	 => data_sig,
		result	 => result_sig
	);
