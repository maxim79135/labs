or10rez_inst : or10rez PORT MAP (
		data	 => data_sig,
		result	 => result_sig
	);
