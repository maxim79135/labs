xor21_inst : xor21 PORT MAP (
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		result	 => result_sig
	);
