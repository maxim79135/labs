sm1_inst : sm1 PORT MAP (
		cin	 => cin_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
